-------------------------------------------------------------------------------
-- File       : AppDataProcessor.vhd
-- Company    : SLAC National Accelerator Laboratory
-------------------------------------------------------------------------------
-- Description: AppDataProcessor File
-------------------------------------------------------------------------------
-- This file is part of 'axi-pcie-core'.
-- It is subject to the license terms in the LICENSE.txt file found in the 
-- top-level directory of this distribution and at: 
--    https://confluence.slac.stanford.edu/display/ppareg/LICENSE.html. 
-- No part of 'axi-pcie-core', including this file, 
-- may be copied, modified, propagated, or distributed except according to 
-- the terms contained in the LICENSE.txt file.
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

use work.StdRtlPkg.all;

use work.AxiPkg.all;
use work.AxiLitePkg.all;
use work.AxiStreamPkg.all;
use work.AppPkg.all;

library unisim;
use unisim.vcomponents.all;

entity AppDataProcessor is
   generic (
      TPD_G            : time             := 1 ns;
      SW_LOOPBACK_G    : boolean          := false;
      AXI_BASE_ADDR_G  : slv(31 downto 0));
   port (
      -- -- Streaming Interfaces
      linkUp          : in  sl;
      sAxisMaster     : in  AxiStreamMasterType;
      sAxisSlave      : out AxiStreamSlaveType;
      mAxisMaster     : out AxiStreamMasterType;
      mAxisSlave      : in  AxiStreamSlaveType;
      loopbackMaster  : in  AxiStreamMasterType;
      loopbackSlave   : out AxiStreamSlaveType;
      -- AXI-Lite Interface
      axilClk         : in  sl;
      axilRst         : in  sl;
      axilReadMaster  : in  AxiLiteReadMasterType;
      axilReadSlave   : out AxiLiteReadSlaveType;
      axilWriteMaster : in  AxiLiteWriteMasterType;
      axilWriteSlave  : out AxiLiteWriteSlaveType);
end AppDataProcessor;

architecture mapping of AppDataProcessor is

begin

   ------------------------------
   -- Placeholder for future code
   ------------------------------
   SW_LOOPBACK : if SW_LOOPBACK_G generate

      mAxisMaster    <= loopbackMaster;
      sAxisSlave     <= AXI_STREAM_SLAVE_FORCE_C;
      loopbackSlave  <= mAxisSlave;

   end generate;

   FW_LOOPBACK : if (not SW_LOOPBACK_G) generate

      mAxisMaster    <= sAxisMaster;
      sAxisSlave     <= mAxisSlave;
      loopbackSlave  <= AXI_STREAM_SLAVE_FORCE_C;

   end generate;

   axilReadSlave  <= AXI_LITE_READ_SLAVE_EMPTY_DECERR_C;
   axilWriteSlave <= AXI_LITE_WRITE_SLAVE_EMPTY_DECERR_C;

end mapping;
